`ifndef _range_sensor_map_svh
`define _range_sensor_map_svh
   
`define SYS_CLK_FREQ 100

`define BRIDGE_BASE 0xc0000000

`define S0_RANGE_SENSOR 0
`define S1_RANGE_SENSOR 1
`define S2_RANGE_SENSOR 2
`define S3_RANGE_SENSOR 3

`endif